-- lab2.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity lab2_top is
	port (
		clk                          : in  std_logic                    := '0'; --                       clk.clk
		seg : out std_logic_vector(6 downto 0);        -- pio_0_external_connection.export
		seg1 : out std_logic_vector(6 downto 0);
		seg2 : out std_logic_vector(6 downto 0);
		reset                   : in  std_logic                    := '0'  --                     reset.reset_n
	);
end entity lab2_top;


architecture arch of lab2_top is
	component Exo2_ESN_sys is
		port (
			clk_clk                          : in  std_logic                    := 'X'; -- clk
			reset_reset_n                    : in  std_logic                    := 'X'; -- reset_n
			pio_0_external_connection_export : out std_logic_vector(3 downto 0);         -- export
			pio_1_external_connection_export : out std_logic_vector(3 downto 0);         -- export
		   pio_2_external_connection_export : out std_logic_vector(3 downto 0)
		);
	end component Exo2_ESN_sys;
	
	component BCD7SEG is
		 port (
			bin_in : in  STD_LOGIC_VECTOR (3 downto 0);
			seg_out : out  STD_LOGIC_VECTOR (6 downto 0));
	end component BCD7SEG;


signal s0 : std_logic_vector(3 downto 0);
signal s1 : std_logic_vector(3 downto 0);
signal s2 : std_logic_vector(3 downto 0);
begin
	u0 : component Exo2_ESN_sys
		port map (
			clk_clk                          => clk,                          --                       clk.clk
			reset_reset_n                    => reset,                    --                     reset.reset_n
			pio_0_external_connection_export => s0,  -- pio_0_external_connection.export
		   pio_1_external_connection_export => s1,
			pio_2_external_connection_export => s2
		);
		
	u1 : component BCD7SEG
		port map (
			bin_in                     => s0,  
			seg_out                    => seg
		);

	u2 : component BCD7SEG
		port map (
			bin_in                     => s1,  
			seg_out                    => seg1
		);
		
	u3 : component BCD7SEG
		port map (
			bin_in                     => s2,  
			seg_out                    => seg2
		);
	end architecture arch;